
    /* verilator lint_off WIDTH */
    /* verilator lint_off CASEINCOMPLETE */
    `include "bsg_defines.v"
    `include "../bsg_misc/bsg_idiv_iterative.v"
    `include "../bsg_misc/bsg_dff_en.v"
    `include "../bsg_misc/bsg_mux_one_hot.v"
    `include "../bsg_misc/bsg_adder_cin.v"
    `include "../bsg_misc/bsg_idiv_iterative_controller.v"
    `include "../bsg_misc/bsg_counter_clear_up.v"
    /* verilator lint_on WIDTH */
    /* verilator lint_on CASEINCOMPLETE */

    module bsg_tanh #(parameter neg_prec_p=6, posi_prec_p=12, extr_iter_p=1, ans_width_p = 32, ang_width_p = 21, precision=16)
    (
    input clk_i
    ,input signed [ang_width_p-1:0] ang_i
    ,input ready_i
    ,input val_i
    ,input reset_i
    ,output signed [ans_width_p-1:0] tanh_o
    ,output ready_o
    ,output val_o
    );

    logic signed [ans_width_p-1:0] sinh, cosh, tanh_r, tanh_n;
    logic sincosReady, sincosDone, tanReady, tanDone, sincos_val_i, tan_val_i, bypass;
    
    
  
    /* state logic */
    enum logic [1:0] {eWAIT, eBUSY1, eBUSY2, eDONE} state_r, state_n;

    always_comb begin
        state_n = state_r;
        case (state_r)
            eWAIT: begin
                if (ready_o && val_i) begin 
                    if (bypass) state_n = eDONE;
                    else        state_n = eBUSY1;
                end
            end
            eBUSY1: begin
                if (bypass) state_n = eDONE;
                else if (sincosDone && tanReady) state_n = eBUSY2;
            end
            eBUSY2: begin
                if (bypass || tanDone) state_n = eDONE;
            end
            eDONE: begin
                if (ready_i) state_n = eWAIT;
            end
            default: state_n = eWAIT;
        endcase
    end

    always_ff @(posedge clk_i) begin
        state_r <= state_n;
    end

    /* bypass if tanh ~= 1 */
    assign bypass = (ang_i > { {(ang_width_p-precision-2){1'b0}}, 5'b11111, {(precision-3){1'b0}} });
    assign sincos_val_i = val_i && ~bypass;
    assign tan_val_i = (sincosDone && (state_r == eBUSY1)) && ~bypass;

    /* sinh cosh module */
    bsg_cordic_sine_cosine_hyperbolic #(.neg_prec_p, .posi_prec_p, .extr_iter_p, .ans_width_p, .ang_width_p) sinhcosh
    (
     .clk_i
    ,.ang_i
    ,.ready_i   (tanReady && (state_r == eWAIT))
    ,.val_i     (sincos_val_i)
    ,.sinh_o    (sinh)
    ,.cosh_o    (cosh)
    ,.ready_o   (sincosReady)
    ,.val_o     (sincosDone)
    );

    /* tan divider unit */
    parameter SHFT_AMT = 16;
    logic [ans_width_p+SHFT_AMT-1:0] sinh_shifted, tanh_shifted, remainder_o, tanh_crop; //L shift by 16
    assign sinh_shifted = {SHFT_AMT'('d0), sinh} << SHFT_AMT;

    bsg_idiv_iterative #(.width_p(ans_width_p+SHFT_AMT)) divider
    (
     .clk_i
    ,.reset_i       

    ,.v_i           (tan_val_i)
    ,.ready_and_o   (tanReady) 

    ,.dividend_i    (sinh_shifted)
    ,.divisor_i     ({SHFT_AMT'('d0), cosh})
    ,.signed_div_i  (1)

    ,.v_o           (tanDone)
    ,.quotient_o    (tanh_shifted)
    ,.remainder_o   
    ,.yumi_i        (ready_i)
    );

    /* outbound signals */
    always_comb begin
        //if value of output exceeds 1 (decimal) then hard set to 1, otherwise keep normal output
        if (tanh_shifted[SHFT_AMT] == 1 || bypass)    tanh_n = {{ans_width_p-SHFT_AMT-1{1'b0}}, 1'b1, {SHFT_AMT{1'b0}}};
        else                                tanh_n = tanh_shifted[ans_width_p-1:0];
    end
    //assign tanh_n = tanh_shifted[ans_width_p-1:0];
    assign val_o = state_r == eDONE;
    assign ready_o = (state_r == eWAIT) && (sincosReady);

    always_ff @(posedge clk_i) begin
        if (tanDone || bypass)    tanh_r <= tanh_n;
        else                      tanh_r <= tanh_r;
    end

    assign tanh_o = tanh_r;

    
    endmodule
